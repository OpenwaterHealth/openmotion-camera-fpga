/*
This demo is for the MachXO3-1300E on Lattice Semiconductor Master Link Board.
*/
module top(pin,reset,debug);

output reg [3:0] pin; 	//LEDs
input reset;			// Reset switch
wire clk_hs;
output wire [3:0] debug;

wire clk_osc;			// Signal from internal oscillator i.e ~6.05 MHz
reg [25:0] clk_f = 0; 		//Count Register i.e 2.885 Hz which is visible to human eyes

//------------------------- Internal Oscillator----------------------
// defparam OSCH_inst.NOM_FREQ = "2.08";	// The default frequency is 2.08 MHz
defparam OSCH_inst.NOM_FREQ = "12.09"; 		// Output frequency if internal oscillator will be ~53.2 MHz
OSCH OSCH_inst( 
.STDBY(1'b0), 	// 0=Enabled, 1=Disabled (Standby – Power down oscillator)
.OSC(clk_osc), 	// Output of internal oscillator
.SEDSTDBY()); 	// This signal is not required if not using SED
//-------------------------------------------------------------------


xclk __ (.CLKI(clk_osc), .CLKOP(clk_hs));

//------------------------- Counter----------------------------------
/* 	A counter is used to slow down the clock for LED shifting logic.
	This actually works as a clock divider with a larger value.
	This is needed because the toggling of an LED at 6.05 MHz (165.28 ns) cannot be seen by human eyes.
*/
always @ (posedge clk_osc)
	begin
		clk_f<=clk_f+1'b1;	// Counter
	end
//-------------------------------------------------------------------


	
//------------------------- Shift register --------------------------
/*
	A walking 1s pattern is generated by shifting "1101" left in each clock cycle.
	A synchronous reset is used to bring back the LEDs to initial state.
	The clock to this logic is the 20th bit of the counter register.
	The clock to this logic is a slower clock made using a counter.
*/
	always @ (posedge clk_f[20])	// Frequency of clk_f[20] will be 2.885 Hz
		begin
			if (reset==0)
				pin<="1101"; 		// Initial value of LEDs.
			else 
				pin<={pin[0],pin[3:1]}; // Shifting the LED values to make a walking 1s pattern
		end	
//-------------------------------------------------------------------
wire reset_n_HFCLKOUT;
wire clk_uart;
wire uart;

//	Reset Bridge for clk_osc
reset_bridge rst_brg_osc(
  .clk_i			(clk_hs),// Destination clock
  .ext_resetn_i		( reset ),// Asynchronous reset signal
  .sync_resetn_out	(reset_n_HFCLKOUT)// Synchronized reset signal
);

wire [9:0] test_pixel;
wire test_lv, test_fv;
grayscale_color_bar gs_i(
	.clk        (clk_hs),            // 133.00 MHz clock
    .reset_n    (reset_n_HFCLKOUT),        // Active low reset
    .pixel_out  (test_pixel),// 10-bit grayscale pixel
    .line_valid (test_lv),     // Line valid signal
    .frame_valid(test_fv)     // Frame valid signal
);

wire spi_clk;

wire [9:0] test_pixel_x;
wire test_lv_x, test_fv_x;

signal_buffer lv_buf(clk_hs, ~reset_n_HFCLKOUT, test_lv, test_lv_x);
signal_buffer fv_buf(clk_hs, ~reset_n_HFCLKOUT, test_fv, test_fv_x);
signal_buffer_10 px_buf(clk_hs, ~reset_n_HFCLKOUT, test_pixel, test_pixel_x);


histogram_module histogram_module_i(
	.clk 		(clk_hs),
	.reset		(~reset_n_HFCLKOUT),
	.pixel_data (test_pixel_x),//test_pixel),
	.frame_valid (test_fv_x),//test_fv),
	.line_valid (test_lv_x),//test_lv),
	.spi_clk_i 	(clk_hs),
	.spi_mosi_o (uart),
	.spi_clk_o (spi_clk),
	.debug		(debug)
//	.debug2		(sldata_o)
); 



endmodule